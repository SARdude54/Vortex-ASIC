`timescale 1ps/1ps

module main (
    input logic A,
    output logic B
);

assign B = A;
    
endmodule

